`ifndef __JVS_PKG_SV__
 `define __JVS_PKG_SV__
`include "jvs_defines.sv"

package jvs_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
`include "jvs_files.sv"
endpackage

`endif