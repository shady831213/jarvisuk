`ifndef __JVS_INTERFACES_SV__
 `define __JVS_INTERFACES_SV__
`include "jvs_irq_interfaces.sv"
`endif