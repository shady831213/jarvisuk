`ifndef __JVS_CLK_RST_GROUP_DEFINES_SV__
 `define __JVS_CLK_RST_GROUP_DEFINES_SV__
 `ifndef JVS_MAX_CLK_GROUP_CLK_NUM
  `define JVS_MAX_CLK_GROUP_CLK_NUM 16
 `endif
`endif