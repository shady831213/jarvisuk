`ifndef __JVS_INTERFACES_SV__
 `define __JVS_INTERFACES_SV__
`include "jvs_irq_interfaces.sv"
`include "jvs_clk_rst_group_interfaces.sv"
`endif