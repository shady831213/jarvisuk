`ifndef __JVS_COMMON_FILES_SV__
 `define __JVS_COMMON_FILES_SV__
`include "jvs_common_attr.sv"
`include "jvs_common_type_queue.sv"
`include "jvs_common_condition.sv"
`endif