`ifndef __JVS_IRQ_FILES_SV__
 `define __JVS_IRQ_FILES_SV__
 `include "jvs_irq_trans.sv"
 `include "jvs_msi_monitor.sv"
 `include "jvs_int_monitor.sv"
 `include "jvs_int_driver.sv"
 `include "jvs_int_agent.sv"
 `include "jvs_irq_handler.sv"
 `include "jvs_irq_vir_sequencer.sv"
 `include "jvs_irq_vir_seq.sv"
 `include "jvs_irq_env.sv"
`endif