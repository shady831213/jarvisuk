`ifndef __JVS_CLK_RST_GROUP_INTERFACES_SV__
 `define __JVS_CLK_RST_GROUP_INTERFACES_SV__
`include "jvs_clk_ifs.sv"
`endif