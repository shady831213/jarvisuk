`ifndef __JVS_REGISTER_REGION_TB_SV__
 `define __JVS_REGISTER_REGION_TB_SV__
`include "uvm_macros.svh"
import uvm_pkg::*;
import jvs_pkg::*;


module jvs_register_region_tb();
   initial begin
      run_test();
    end
endmodule

`endif