`ifndef __JVS_CLK_RST_GROUP_FILES_SV__
 `define __JVS_CLK_RST_GROUP_FILES_SV__
 `include "jvs_clk_rst_trans.sv"
 `include "jvs_clk_driver.sv"
 `include "jvs_clk_vir_seqr.sv"
 `include "jvs_clk_agent.sv"
 `include "jvs_clk_env.sv"
`endif