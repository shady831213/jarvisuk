`ifndef __JVS_FILES_SV__
 `define __JVS_FILES_SV__
 `include "jvs_common_files.sv"
 `include "jvs_memory_files.sv"
 `include "jvs_irq_files.sv"
 `include "jvs_register_region_files.sv"
 `include "jvs_clk_rst_group_files.sv"
`endif