`ifndef __JVS_MEMORY_FILES_SV__
 `define __JVS_MEMORY_FILES_SV__
`include "jvs_memory_types.sv"
`include "jvs_memory_model.sv"
`include "jvs_memory_allocator.sv"
`include "jvs_memory_block.sv"
`endif