`ifndef __JVS_REGISTER_REGION_FILES_SV__
 `define __JVS_REGISTER_REGION_FILES_SV__
`include "jvs_reg_resource_manager.sv"
`include "jvs_reg_tree.sv"
`include "jvs_reg_block_wrapper.sv"
`include "jvs_reg_region.sv"
`include "jvs_reg_region_builder.sv"
`include "jvs_reg_region_mapper.sv"
`endif