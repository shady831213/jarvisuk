`ifndef __JVS_IRQ_INTERFACES_SV__
 `define __JVS_IRQ_INTERFACES_SV__
 `include "jvs_int_if.sv"
`endif